`define	MOV_AR      8'b1
`define	MOV_RR_LOAD 8'b10
`define	MOV_RA      8'b11
`define	ADD         8'b10000
`define	SUB         8'b10001
`define	AND         8'b10010
`define	OR          8'b10011
`define	NOT         8'b10100
`define	XOR         8'b10101
`define	RAND        8'b10110
`define	ROR         8'b10111
`define	RXOR        8'b11000
`define	LSL         8'b11001
`define	LSR         8'b11010
`define	ASL         8'b11011
`define	ASR         8'b11100
`define	CSL         8'b11101
`define	CSR         8'b11110
`define	INC         8'b11111
`define	DEC         8'b100000
`define	PUSH        8'b1010000
`define	POP         8'b1010001
`define	SAVEPC      8'b10000000
`define	RECOPC      8'b10000000
